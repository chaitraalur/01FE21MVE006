class  generator
rand transaction trans;
mailbox gen2driver;
initial count();
event ended();
function mailbox=new();
end class
